library verilog;
use verilog.vl_types.all;
entity MaquinaDestadosV1_vlg_vec_tst is
end MaquinaDestadosV1_vlg_vec_tst;
